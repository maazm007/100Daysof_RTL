module Nine_Bit_MUX(Mux_Out,A,B,Sel,Reset);
	input [8:0] A;
	input [8:0] B;
	input Sel, Reset;
	output [8:0] Mux_Out;
	wire w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15;
	assign A[8] = 1'b0;
	and n1(w1,~Sel,A[0]);
	and n2(w2,Sel,B[0]);
	or o1(Mux_Out[0],w1,w2);
	and n3(w3,~Sel,A[1]);
	and n4(w4,Sel,B[1]);
	or o2(Mux_Out[1],w3,w4);
	and n5(w5,~Sel,A[2]);
	and n6(w6,Sel,B[2]);
	or o3(Mux_Out[2],w5,w6);
	and n7(w7,~Sel,A[3]);
	and n8(w8,Sel,B[3]);
	or o4(Mux_Out[3],w7,w8);
	and n9(w9,~Sel,A[4]);
	and n10(w10,Sel,B[4]);
	or o5(Mux_Out[4],w9,w10);
	and n11(w11,~Sel,A[5]);
	and n12(w12,Sel,B[5]);
	or o6(Mux_Out[5],w11,w12);
	and n13(w13,~Sel,A[6]);
	and n14(w14,Sel,B[6]);
	or o7(Mux_Out[6],w13,w14);
	and n15(w15,~Sel,A[7]);
	and n16(w16,Sel,B[7]);
	or o8(Mux_Out[7],w15,w16);
	and n17(w17,~Sel,A[8]);
	and n18(w18,Sel,B[8]);
	or o9(Mux_Out[8],w17,w18);
endmodule
